library verilog;
use verilog.vl_types.all;
entity kamal_lab1_3to8Decoder_vlg_vec_tst is
end kamal_lab1_3to8Decoder_vlg_vec_tst;
