library verilog;
use verilog.vl_types.all;
entity kamal_lab1_8to3Encoder_vlg_sample_tst is
    port(
        kamal_input0    : in     vl_logic;
        kamal_input1    : in     vl_logic;
        kamal_input2    : in     vl_logic;
        kamal_input3    : in     vl_logic;
        kamal_input4    : in     vl_logic;
        kamal_input5    : in     vl_logic;
        kamal_input6    : in     vl_logic;
        kamal_input7    : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end kamal_lab1_8to3Encoder_vlg_sample_tst;
