library verilog;
use verilog.vl_types.all;
entity kamal_lab1_AdderLPM_vlg_sample_tst is
    port(
        dataa           : in     vl_logic_vector(0 downto 0);
        datab           : in     vl_logic_vector(0 downto 0);
        sampler_tx      : out    vl_logic
    );
end kamal_lab1_AdderLPM_vlg_sample_tst;
