library verilog;
use verilog.vl_types.all;
entity kamal_muxLPM_vlg_check_tst is
    port(
        result          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_muxLPM_vlg_check_tst;
