library verilog;
use verilog.vl_types.all;
entity kamal_lab1_3to8Decoder_vlg_check_tst is
    port(
        kamal_outputz0  : in     vl_logic;
        kamal_outputz1  : in     vl_logic;
        kamal_outputz2  : in     vl_logic;
        kamal_outputz3  : in     vl_logic;
        kamal_outputz4  : in     vl_logic;
        kamal_outputz5  : in     vl_logic;
        kamal_outputz6  : in     vl_logic;
        kamal_outputz7  : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_lab1_3to8Decoder_vlg_check_tst;
