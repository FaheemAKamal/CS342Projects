library verilog;
use verilog.vl_types.all;
entity kamal_Lab1_Decoder_vlg_vec_tst is
end kamal_Lab1_Decoder_vlg_vec_tst;
