library verilog;
use verilog.vl_types.all;
entity kamal_lab1_fulladderlpm_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        result          : in     vl_logic_vector(0 downto 0);
        sampler_rx      : in     vl_logic
    );
end kamal_lab1_fulladderlpm_vlg_check_tst;
