library verilog;
use verilog.vl_types.all;
entity kamal_lab1fulladder_vlg_check_tst is
    port(
        kamal_outputCout: in     vl_logic;
        kamal_outputs   : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_lab1fulladder_vlg_check_tst;
