library verilog;
use verilog.vl_types.all;
entity kamal_mux2to1_vlg_vec_tst is
end kamal_mux2to1_vlg_vec_tst;
