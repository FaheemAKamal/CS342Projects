library verilog;
use verilog.vl_types.all;
entity kamal_lab1halfadder is
    port(
        kamal_outputc   : out    vl_logic;
        kamal_inputa    : in     vl_logic;
        kamal_inputb    : in     vl_logic;
        kamal_outputd   : out    vl_logic
    );
end kamal_lab1halfadder;
