library verilog;
use verilog.vl_types.all;
entity kamal_lab1halfadder_vlg_check_tst is
    port(
        kamal_outputc   : in     vl_logic;
        kamal_outputd   : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_lab1halfadder_vlg_check_tst;
