library verilog;
use verilog.vl_types.all;
entity kamal_mux2to1_vlg_check_tst is
    port(
        kamal_outputm   : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_mux2to1_vlg_check_tst;
