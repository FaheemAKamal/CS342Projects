library verilog;
use verilog.vl_types.all;
entity kamal_simpleCircuit_vlg_vec_tst is
end kamal_simpleCircuit_vlg_vec_tst;
