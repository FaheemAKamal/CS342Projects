library verilog;
use verilog.vl_types.all;
entity kamal_simpleCircuit_vlg_check_tst is
    port(
        kamal_outputf   : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_simpleCircuit_vlg_check_tst;
