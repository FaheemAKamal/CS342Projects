library verilog;
use verilog.vl_types.all;
entity kamal_muxLPM_vlg_vec_tst is
end kamal_muxLPM_vlg_vec_tst;
