library verilog;
use verilog.vl_types.all;
entity kamal_lab1_8to3Encoder_vlg_vec_tst is
end kamal_lab1_8to3Encoder_vlg_vec_tst;
