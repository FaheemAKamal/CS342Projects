library verilog;
use verilog.vl_types.all;
entity kamal_lab1_3to8Decoder_vlg_sample_tst is
    port(
        kamal_input1    : in     vl_logic;
        kamal_input2    : in     vl_logic;
        kamal_input3    : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end kamal_lab1_3to8Decoder_vlg_sample_tst;
