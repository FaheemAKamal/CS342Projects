library verilog;
use verilog.vl_types.all;
entity kamal_Lab1_Decoder_vlg_check_tst is
    port(
        eq7             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_Lab1_Decoder_vlg_check_tst;
