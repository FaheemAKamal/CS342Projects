library verilog;
use verilog.vl_types.all;
entity kamal_lab1_8to3Encoder_vlg_check_tst is
    port(
        kamal_outputY1  : in     vl_logic;
        kamal_outputY2  : in     vl_logic;
        kamal_outputY3  : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end kamal_lab1_8to3Encoder_vlg_check_tst;
