library verilog;
use verilog.vl_types.all;
entity kamal_lab1_8to3Encoder is
    port(
        kamal_outputY1  : out    vl_logic;
        kamal_input4    : in     vl_logic;
        kamal_input6    : in     vl_logic;
        kamal_input7    : in     vl_logic;
        kamal_input5    : in     vl_logic;
        kamal_outputY2  : out    vl_logic;
        kamal_input2    : in     vl_logic;
        kamal_input3    : in     vl_logic;
        kamal_outputY3  : out    vl_logic;
        kamal_input1    : in     vl_logic;
        kamal_input0    : in     vl_logic
    );
end kamal_lab1_8to3Encoder;
