library verilog;
use verilog.vl_types.all;
entity kamal_lab1_3to8Decoder is
    port(
        kamal_outputz0  : out    vl_logic;
        kamal_input1    : in     vl_logic;
        kamal_input2    : in     vl_logic;
        kamal_input3    : in     vl_logic;
        kamal_outputz1  : out    vl_logic;
        kamal_outputz2  : out    vl_logic;
        kamal_outputz3  : out    vl_logic;
        kamal_outputz4  : out    vl_logic;
        kamal_outputz5  : out    vl_logic;
        kamal_outputz6  : out    vl_logic;
        kamal_outputz7  : out    vl_logic
    );
end kamal_lab1_3to8Decoder;
